netcdf argo-trajectory-v2.1-spec {

//@ DATA_TYPE = "Argo trajectory"
//@ FORMAT_VERSION   = "2.2"
//@ HANDBOOK_VERSION = "1.2"
//@ REFERENCE_DATE_TIME = "19500101000000"
//@ $Revision: 657 $
//@ $Date: 2017-04-24 16:48:54 +0000 (Mon, 24 Apr 2017) $

dimensions:
	DATE_TIME = 14;
	STRING256 = 256;
	STRING64 = 64;
	STRING32 = 32;
	STRING16 = 16;
	STRING8 = 8;
	STRING4 = 4;
	STRING2 = 2;

	N_PARAM = _unspecified_;
	N_CYCLE = _unspecified_;
	N_HISTORY = _unspecified_;
	N_MEASUREMENT = UNLIMITED;

variables:
	char DATA_TYPE(STRING16);
		DATA_TYPE:long_name = "Data type";
		DATA_TYPE:_FillValue = " ";
	char FORMAT_VERSION(STRING4);
		FORMAT_VERSION:long_name = "File format version";
		FORMAT_VERSION:_FillValue = " ";
	char HANDBOOK_VERSION(STRING4);
		HANDBOOK_VERSION:long_name = "Data handbook version";
		HANDBOOK_VERSION:_FillValue = " ";
	char REFERENCE_DATE_TIME(DATE_TIME);
		REFERENCE_DATE_TIME:long_name = "Date of reference for Julian days";
		REFERENCE_DATE_TIME:conventions = "YYYYMMDDHHMISS";
		REFERENCE_DATE_TIME:_FillValue = " ";
	char DATE_CREATION(DATE_TIME);
		DATE_CREATION:long_name = "Date of file creation";
		DATE_CREATION:conventions = "YYYYMMDDHHMISS";
		DATE_CREATION:_FillValue = " ";
	char DATE_UPDATE(DATE_TIME);
		DATE_UPDATE:long_name = "Date of update of this file";
		DATE_UPDATE:conventions = "YYYYMMDDHHMISS";
		DATE_UPDATE:_FillValue = " ";
	char PLATFORM_NUMBER(STRING8);
		PLATFORM_NUMBER:long_name = "Float unique identifier";
		PLATFORM_NUMBER:conventions = "WMO float identifier : A9IIIII";
		PLATFORM_NUMBER:_FillValue = " ";
	char PROJECT_NAME(STRING64);
		PROJECT_NAME:long_name = "Name of the project";
		PROJECT_NAME:_FillValue = " ";
	char PI_NAME (STRING64);
		PI_NAME:long_name = "Name of the principal investigator";
		PI_NAME:_FillValue = " ";
	char TRAJECTORY_PARAMETERS(N_PARAM, STRING16);
		TRAJECTORY_PARAMETERS:long_name = "List of available parameters for the station";
		TRAJECTORY_PARAMETERS:conventions = "Argo reference table 3";
		TRAJECTORY_PARAMETERS:_FillValue = " ";
	char DATA_CENTRE(STRING2);
		DATA_CENTRE:long_name = "Data centre in charge of float data processing";
		DATA_CENTRE:conventions = "Argo reference table 4";
		DATA_CENTRE:_FillValue = " ";
	char DATA_STATE_INDICATOR(STRING4);
		DATA_STATE_INDICATOR:long_name = "Degree of processing the data have passed through";
		DATA_STATE_INDICATOR:conventions = "Argo reference table 6";
		DATA_STATE_INDICATOR:_FillValue = " ";
	char INST_REFERENCE(STRING64);
		INST_REFERENCE:long_name = "Instrument type";
		INST_REFERENCE:conventions = "Brand, type, serial number";
		INST_REFERENCE:_FillValue = " ";
	char WMO_INST_TYPE(STRING4);
		WMO_INST_TYPE:long_name = "Coded instrument type";
		WMO_INST_TYPE:conventions = "Argo reference table 8";
		WMO_INST_TYPE:_FillValue = " ";
	char POSITIONING_SYSTEM(STRING8);
		POSITIONING_SYSTEM:long_name = "Positioning system";
		POSITIONING_SYSTEM:_FillValue = " ";
	double JULD(N_MEASUREMENT);
		JULD:long_name = "Julian day (UTC) of each measurement relative to REFERENCE_DATE_TIME";
                JULD:standard_name = "time" ; 
		JULD:units = "days since 1950-01-01 00:00:00 UTC";
		JULD:conventions = "Relative julian days with decimal part (as parts of the day)";
		JULD:_FillValue = 999999.;
                JULD:axis = "T" ; 
	char JULD_QC(N_MEASUREMENT);
		JULD_QC:long_name = "Quality on date and time";
		JULD_QC:conventions = "Argo reference table 2";
		JULD_QC:_FillValue = " ";
	double LATITUDE(N_MEASUREMENT);
		LATITUDE:long_name = "Latitude of each location";
                LATITUDE:standard_name = "latitude"; 
		LATITUDE:units = "degree_north";
		LATITUDE:_FillValue = 99999.;
		LATITUDE:valid_min = -90.;
		LATITUDE:valid_max = 90.;
                LATITUDE:axis = "Y" ;
	double LONGITUDE(N_MEASUREMENT);
		LONGITUDE:long_name = "Longitude of each location";
                LONGITUDE:standard_name = "longitude" ;
		LONGITUDE:units = "degree_east";
		LONGITUDE:_FillValue = 99999.;
		LONGITUDE:valid_min = -180.;
		LONGITUDE:valid_max = 180.;
                LONGITUDE:axis = "X" ;
	char POSITION_ACCURACY(N_MEASUREMENT);
		POSITION_ACCURACY:long_name = "Estimated accuracy in latitude and longitude";
		POSITION_ACCURACY:conventions = "Argo reference table 5";
		POSITION_ACCURACY:_FillValue = " ";
	char POSITION_QC(N_MEASUREMENT);
		POSITION_QC:long_name = "Quality on position";
		POSITION_QC:conventions = "Argo reference table 2";
		POSITION_QC:_FillValue = " ";
	int CYCLE_NUMBER(N_MEASUREMENT);
		CYCLE_NUMBER:long_name = "Float cycle number of the measurement";
		CYCLE_NUMBER:conventions = "0..N, 0 : launch cycle, 1 : first complete cycle";
		CYCLE_NUMBER:_FillValue = 99999;
	int MEASUREMENT_CODE (N_MEASUREMENT);
		MEASUREMENT_CODE:long_name = "Code referring to a measurement event in the cycle";
		MEASUREMENT_CODE:conventions = "Argo reference table 15";
		MEASUREMENT_CODE:_FillValue = 99999;

// Physical parameters added via argo-physical_params*

	double JULD_ASCENT_START(N_CYCLE);
		JULD_ASCENT_START:long_name = "Start date of the ascending profile";
		JULD_ASCENT_START:units = "days since 1950-01-01 00:00:00 UTC";
		JULD_ASCENT_START:conventions = "Relative julian days with decimal part (as part of day)";
		JULD_ASCENT_START:_FillValue = 999999.;
	char JULD_ASCENT_START_STATUS(N_CYCLE);
		JULD_ASCENT_START_STATUS:conventions = "0 : Nominal, 1 : Estimated, 2 : Transmitted";
		JULD_ASCENT_START_STATUS:_FillValue = " ";
	double JULD_ASCENT_END(N_CYCLE);
		JULD_ASCENT_END:long_name = "End date of the ascending profile";
		JULD_ASCENT_END:units = "days since 1950-01-01 00:00:00 UTC";
		JULD_ASCENT_END:conventions = "Relative julian days with decimal part (as part of day)";
		JULD_ASCENT_END:_FillValue = 999999.;
	char JULD_ASCENT_END_STATUS(N_CYCLE);
		JULD_ASCENT_END_STATUS:conventions = "0 : Nominal, 1 : Estimated, 2 : Transmitted";
		JULD_ASCENT_END_STATUS:_FillValue = " ";
	double JULD_DESCENT_START(N_CYCLE);
		JULD_DESCENT_START:long_name = "Descent start date of the cycle";
		JULD_DESCENT_START:units = "days since 1950-01-01 00:00:00 UTC";
		JULD_DESCENT_START:conventions = "Relative julian days with decimal part (as part of day)";
		JULD_DESCENT_START:_FillValue = 999999.;
	char JULD_DESCENT_START_STATUS(N_CYCLE);
		JULD_DESCENT_START_STATUS:conventions = "0 : Nominal, 1 : Estimated, 2 : Transmitted";
		JULD_DESCENT_START_STATUS:_FillValue = " ";
	double JULD_DESCENT_END(N_CYCLE);
		JULD_DESCENT_END:long_name = "Descent end date of the cycle";
		JULD_DESCENT_END:units = "days since 1950-01-01 00:00:00 UTC";
		JULD_DESCENT_END:conventions = "Relative julian days with decimal part (as part of day)";
		JULD_DESCENT_END:_FillValue = 999999.;
	char JULD_DESCENT_END_STATUS(N_CYCLE);
		JULD_DESCENT_END_STATUS:conventions = "0 : Nominal, 1 : Estimated, 2 : Transmitted";
		JULD_DESCENT_END_STATUS:_FillValue = " ";

	double JULD_TRANSMISSION_START(N_CYCLE);
		JULD_TRANSMISSION_START:long_name = "Start date of transmission";
		JULD_TRANSMISSION_START:units = "days since 1950-01-01 00:00:00 UTC";
		JULD_TRANSMISSION_START:conventions = "Relative julian days with decimal part (as part of day)";
		JULD_TRANSMISSION_START:_FillValue=999999.;
	char JULD_TRANSMISSION_START_STATUS(N_CYCLE);
		JULD_TRANSMISSION_START_STATUS:conventions = "0 : Nominal, 1 : Estimated, 2 : Transmitted";
		JULD_TRANSMISSION_START_STATUS:_FillValue = " ";
	double JULD_FIRST_STABILIZATION(N_CYCLE);
		JULD_FIRST_STABILIZATION:long_name = "Time of float's first stabilization after leaving the surface";
		JULD_FIRST_STABILIZATION:units = "days since 1950-01-01 00:00:00 UTC";
		JULD_FIRST_STABILIZATION:conventions = "Relative julian days with decimal part (as part of day)";
		JULD_FIRST_STABILIZATION:_FillValue=999999.;
	char JULD_FIRST_STABILIZATION_STATUS(N_CYCLE);
		JULD_FIRST_STABILIZATION_STATUS:conventions = "0 : Nominal, 1 : Estimated, 2 : Transmitted";
		JULD_FIRST_STABILIZATION_STATUS:_FillValue = " ";
	double JULD_DEEP_DESCENT_START(N_CYCLE);
		JULD_DEEP_DESCENT_START:long_name = "Deep Descent start date of the cycle";
		JULD_DEEP_DESCENT_START:units = "days since 1950-01-01 00:00:00 UTC";
		JULD_DEEP_DESCENT_START:conventions = "Relative julian days with decimal part (as part of day)";
		JULD_DEEP_DESCENT_START:_FillValue=999999.;
	char JULD_DEEP_DESCENT_START_STATUS(N_CYCLE);
		JULD_DEEP_DESCENT_START_STATUS:conventions = "0 : Nominal, 1 : Estimated, 2 : Transmitted";
		JULD_DEEP_DESCENT_START_STATUS:_FillValue = " ";
	double JULD_DEEP_DESCENT_END(N_CYCLE);
		JULD_DEEP_DESCENT_END:long_name = "Deep Descent end date of the cycle";
		JULD_DEEP_DESCENT_END:units = "days since 1950-01-01 00:00:00 UTC";
		JULD_DEEP_DESCENT_END:conventions = "Relative julian days with decimal part (as part of day)";
		JULD_DEEP_DESCENT_END:_FillValue=999999.;
	char JULD_DEEP_DESCENT_END_STATUS(N_CYCLE);
		JULD_DEEP_DESCENT_END_STATUS:conventions = "0 : Nominal, 1 : Estimated, 2 : Transmitted";
		JULD_DEEP_DESCENT_END_STATUS:_FillValue = " ";
	double JULD_TRANSMISSION_END(N_CYCLE);
		JULD_TRANSMISSION_END:long_name = "Transmission end date";
		JULD_TRANSMISSION_END:units = "days since 1950-01-01 00:00:00 UTC";
		JULD_TRANSMISSION_END:conventions = "Relative julian days with decimal part (as part of day)";
		JULD_TRANSMISSION_END:_FillValue=999999.;
	char JULD_TRANSMISSION_END_STATUS(N_CYCLE);
		JULD_TRANSMISSION_END_STATUS:conventions = "0 : Nominal, 1 : Estimated, 2 : Transmitted";
		JULD_TRANSMISSION_END_STATUS:_FillValue = " ";
	char GROUNDED(N_CYCLE);
		GROUNDED:long_name = "Did the profiler touch the ground for that cycle";
                GROUNDED:conventions = "Y,P,N,U";
		GROUNDED:_FillValue = " ";
	int CONFIG_MISSION_NUMBER (N_CYCLE);
		CONFIG_MISSION_NUMBER:long_name = "mission number of unique cycles performed by the float";
		CONFIG_MISSION_NUMBER:_FillValue = 99999;
	int CYCLE_NUMBER_ACTUAL(N_CYCLE);
		CYCLE_NUMBER_ACTUAL:long_name = "Float cycle number of the measurement";
		CYCLE_NUMBER_ACTUAL:conventions = "0...N, 0 : lauch cycle, 1 : first complete cycle";
		CYCLE_NUMBER_ACTUAL:_FillValue = 99999;
	char DATA_MODE(N_CYCLE);
		DATA_MODE:long_name = "Delayed mode or real time data";
		DATA_MODE:conventions = "R : real time; D : delayed mode; A : real time with adjustment";
		DATA_MODE:_FillValue = " ";

	char HISTORY_INSTITUTION (N_HISTORY, STRING4);
		HISTORY_INSTITUTION:long_name = "Institution which performed action";
		HISTORY_INSTITUTION:conventions = "Argo reference table 4";
		HISTORY_INSTITUTION:_FillValue = " ";
	char HISTORY_STEP(N_HISTORY, STRING4);
		HISTORY_STEP:long_name = "Step in data processing";
		HISTORY_STEP:conventions = "Argo reference table 12";
		HISTORY_STEP:_FillValue = " ";
	char HISTORY_SOFTWARE(N_HISTORY, STRING4);
		HISTORY_SOFTWARE:long_name = "Name of software which performed action";
		HISTORY_SOFTWARE:conventions = "Institution dependent";
		HISTORY_SOFTWARE:_FillValue = " ";
	char HISTORY_SOFTWARE_RELEASE(N_HISTORY, STRING4);
		HISTORY_SOFTWARE_RELEASE:long_name = "Version/release of software which performed action";
		HISTORY_SOFTWARE_RELEASE:conventions = "Institution dependent";
		HISTORY_SOFTWARE_RELEASE:_FillValue = " ";
	char HISTORY_REFERENCE(N_HISTORY, STRING64);
		HISTORY_REFERENCE:long_name = "Reference of database";
		HISTORY_REFERENCE:conventions = "Institution dependent";
		HISTORY_REFERENCE:_FillValue = " ";
	char HISTORY_DATE(N_HISTORY, DATE_TIME);
		HISTORY_DATE:long_name = "Date the history record was created";
		HISTORY_DATE:conventions = "YYYYMMDDHHMISS";
		HISTORY_DATE:_FillValue = " ";
	char HISTORY_ACTION(N_HISTORY, STRING4);
		HISTORY_ACTION:long_name = "Action performed on data";
		HISTORY_ACTION:conventions = "Argo reference table 7";
		HISTORY_ACTION:_FillValue = " ";
	char HISTORY_PARAMETER(N_HISTORY, STRING16);
		HISTORY_PARAMETER:long_name = "Station parameter action is performed on";
		HISTORY_PARAMETER:conventions = "Argo reference table 3";
		HISTORY_PARAMETER:_FillValue = " ";
	float HISTORY_PREVIOUS_VALUE(N_HISTORY);
		HISTORY_PREVIOUS_VALUE:long_name = "Parameter/Flag previous value before action";
		HISTORY_PREVIOUS_VALUE:_FillValue = 99999.f;
        char HISTORY_INDEX_DIMENSION(N_HISTORY);
	int HISTORY_START_INDEX(N_HISTORY);
		HISTORY_START_INDEX:long_name = "Start index action applied on";
		HISTORY_START_INDEX:_FillValue = 99999;
	int HISTORY_STOP_INDEX(N_HISTORY);
		HISTORY_STOP_INDEX:long_name = "Stop index action applied on";
		HISTORY_STOP_INDEX:_FillValue = 99999;
	char HISTORY_QCTEST(N_HISTORY, STRING16);
		HISTORY_QCTEST:long_name = "Documentation of tests performed, tests failed (in hex form)";
		HISTORY_QCTEST:conventions = "Write tests performed when ACTION=QCP$; tests failed when ACTION=QCF$";
		HISTORY_QCTEST:_FillValue = " ";
}
