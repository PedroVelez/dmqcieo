netcdf argo-technical-v2.1-spec {

//@ DATA_TYPE = "Argo technical"
//@ FORMAT_VERSION   = "2.3"
//@ HANDBOOK_VERSION = "1.2"
//@ $Revision: 657 $
//@ $Date: 2017-04-24 16:48:54 +0000 (Mon, 24 Apr 2017) $

dimensions:

	DATE_TIME = 14;
	STRING128 = 128;
	STRING64 = 64;
	STRING32 = 32;
	STRING16 = 16;
	STRING8 = 8;
	STRING4 = 4;
	STRING2 = 2;
	N_TECH_PARAM = UNLIMITED;

variables:
	char PLATFORM_NUMBER(STRING8);
		PLATFORM_NUMBER:long_name = "Float unique identifier";
		PLATFORM_NUMBER:conventions = "WMO float identifier : A9IIIII";
		PLATFORM_NUMBER:_FillValue = " ";
	char DATA_TYPE(STRING32);
// AB 20120820
//		DATA_TYPE:comment = "Data type";
		DATA_TYPE:_FillValue = " "
	char FORMAT_VERSION(STRING4);
// AB 20120820
//		FORMAT_VERSION:comment = "File format version";
		FORMAT_VERSION:_FillValue = " ";
	char HANDBOOK_VERSION(STRING4);
// AB 20120820
//		HANDBOOK_VERSION:comment = "Data handbook version";
		HANDBOOK_VERSION:_FillValue = " ";
	char DATA_CENTRE(STRING2);
		DATA_CENTRE:long_name = "Data centre in charge of float data processing";
		DATA_CENTRE:conventions = "Argo reference table 4";
		DATA_CENTRE:_FillValue = " ";
	char DATE_CREATION(DATE_TIME);
// AB 20120820
//		DATE_CREATION:comment = "Date of file creation";
		DATE_CREATION:conventions = "YYYYMMDDHHMISS";
		DATE_CREATION:_FillValue = " ";
	char DATE_UPDATE(DATE_TIME);
		DATE_UPDATE:long_name = "Date of update of this file";
		DATE_UPDATE:conventions = "YYYYMMDDHHMISS";
		DATE_UPDATE:_FillValue = " ";
	char TECHNICAL_PARAMETER_NAME(N_TECH_PARAM, STRING128);
		TECHNICAL_PARAMETER_NAME:long_name = "Name of technical parameter";
		TECHNICAL_PARAMETER_NAME:_FillValue = " ";
	char TECHNICAL_PARAMETER_VALUE(N_TECH_PARAM, STRING128);
		TECHNICAL_PARAMETER_VALUE:long_name = "Value of technical parameter";
		TECHNICAL_PARAMETER_VALUE:_FillValue = " ";
	int CYCLE_NUMBER(N_TECH_PARAM);
	        CYCLE_NUMBER:long_name = "Float cycle number";
	        CYCLE_NUMBER:conventions = "0..N, 0 : launch cycle (if exists), 1 : first complete cycle";
		CYCLE_NUMBER:_FillValue = 99999;

}
